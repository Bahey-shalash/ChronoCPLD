--==============================================================================
--== Logisim-evolution goes FPGA automatic generated VHDL code                ==
--== https://github.com/logisim-evolution/                                    ==
--==                                                                          ==
--==                                                                          ==
--== Project   : project_Finale                                               ==
--== Component : NOR_GATE_21_INPUTS                                           ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY NOR_GATE_21_INPUTS IS
   GENERIC ( BubblesMask : std_logic_vector );
   PORT ( input1  : IN  std_logic;
          input10 : IN  std_logic;
          input11 : IN  std_logic;
          input12 : IN  std_logic;
          input13 : IN  std_logic;
          input14 : IN  std_logic;
          input15 : IN  std_logic;
          input16 : IN  std_logic;
          input17 : IN  std_logic;
          input18 : IN  std_logic;
          input19 : IN  std_logic;
          input2  : IN  std_logic;
          input20 : IN  std_logic;
          input21 : IN  std_logic;
          input3  : IN  std_logic;
          input4  : IN  std_logic;
          input5  : IN  std_logic;
          input6  : IN  std_logic;
          input7  : IN  std_logic;
          input8  : IN  std_logic;
          input9  : IN  std_logic;
          result  : OUT std_logic );
END ENTITY NOR_GATE_21_INPUTS;
